
** sch_path: /home/anilk/DC_CHAR/DC_PFET1v8.sch
**.subckt DC_PFET1v8
VSG GND VG 2
XM1 VD VG GND GND sky130_fd_pr__pfet_01v8 L=2 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
VDg VD GND -2


**** begin user architecture code

.lib /usr/local/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt


.save all
.save i(vs)
.save @m.xm1.msky130_fd_pr__pfet_01v8[gm]
.save @m.xm1.msky130_fd_pr__pfet_01v8[id]
.save @m.xm1.msky130_fd_pr__pfet_01v8[vth]
.save @m.xm1.msky130_fd_pr__pfet_01v8[gds]
.save @m.xm1.msky130_fd_pr__pfet_01v8[cgg]
.save @m.xm1.msky130_fd_pr__pfet_01v8[cgs]
.save @m.xm1.msky130_fd_pr__pfet_01v8[cbg]
.save @m.xm1.msky130_fd_pr__pfet_01v8[cdd]
.save @m.xm1.msky130_fd_pr__pfet_01v8[cds]
.save @m.xm1.msky130_fd_pr__pfet_01v8[cgd]
.save @m.xm1.msky130_fd_pr__pfet_01v8[gm]

.option filetype=ascii

.control
    dc VSG 0 2 0.01 VDg -0.1 -1 -0.1
    let gm = @m.xm1.msky130_fd_pr__pfet_01v8[gm]
    let idbyw = @m.xm1.msky130_fd_pr__pfet_01v8[id]/2
    let gmbyid = @m.xm1.msky130_fd_pr__pfet_01v8[gm]/@m.xm1.msky130_fd_pr__pfet_01v8[id]
    let gmbygds = @m.xm1.msky130_fd_pr__pfet_01v8[gm]/@m.xm1.msky130_fd_pr__pfet_01v8[gds]
    let ft = @m.xm1.msky130_fd_pr__pfet_01v8[gm]/@m.xm1.msky130_fd_pr__pfet_01v8[cgg]
    let cgg = @m.xm1.msky130_fd_pr__pfet_01v8[cgg]
    let gds = @m.xm1.msky130_fd_pr__pfet_01v8[gds]
    let Voverdrive = -v(vg)-@m.xm1.msky130_fd_pr__pfet_01v8[vth]
    *let vth = @m.xm1.msky130_fd_pr__pfet_01v8[vth]
    wrdata /home/anilk/SKYWATER130_GMID/PMOS/pmos_data/gmid_pmos_output.txt gm idbyw gmbyid gmbygds ft cgg gds Voverdrive
    *plot idbyw
    quit
.endc

.end
